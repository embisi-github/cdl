/*a Copyright
  
  This file 'hierarchy_test_harness.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/

/*a Includes
 */
include "hierarchy.h"

/*a Constants
 */
constant integer width=16;

/*a Module
 */
module hierarchy_test_harness( clock io_clock,
                               input bit io_reset,
                               input bit[width] vector_input_0,
                               input bit[width] vector_input_1,
                               output bit[width] vector_output_0,
                               output bit[width] vector_output_1 )
    "This module is a wrapper around the hierarchy test modules"
{
    net bit last_value;
    net bit value;
    net bit next_value;
    instances "Instances":
        {
            hierarchy h( int_clock<-io_clock,
                         int_reset<=io_reset,
                         clear<=vector_input_0[0],
                         store<=vector_input_0[1],
                         data<=vector_input_0[2],
                         last_value=>last_value,
                         value=>value,
                         next_value=>next_value );
        }
    drive_outputs "Drive outputs":
        {
            vector_output_1 = 0;
            vector_output_0 = 0;
            vector_output_0[0] = last_value;
            vector_output_0[1] = value;
            vector_output_0[2] = next_value;
        }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

