/*a Copyright
  
  This file 'hierarchy_struct_test_harness.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/

/*a Includes
 */
include "hierarchy_struct.h"

/*a Constants
 */
constant integer width=16;

/*a Module
 */
module hierarchy_struct_test_harness( clock io_clock,
                                      input bit io_reset,
                                      input bit[width] vector_input_0,
                                      input bit[width] vector_input_1,
                                      output bit[width] vector_output_0,
                                      output bit[width] vector_output_1 )
"
This module is a wrapper around the hierarchy test modules

Here is a table of input vectors to result (x=current value)

0 000 -> x
1 001 -> 0
2 010 -> 0
3 011 -> 0
4 100 -> x
5 101 -> 0
6 110 -> 1
7 111 -> 0
"
{
    net t_h_struct out;
    comb t_h_struct in;
    
    instances "Instances":
        {
            in.s.x = vector_input_0[0] ? 1b0 : ( vector_input_0[1]?vector_input_0[2]:out.s.x ); // next_value = clear?0:(store?new:old)
            in.s.y = out.s.x; // last_value
            in.c = out.s.y; // for something
            hierarchy_struct h_s( int_clock<-io_clock,
                                  int_reset<=io_reset,
                                  in <= in,
                                  out => out );
        }
    drive_outputs "Drive outputs":
        {
            vector_output_1 = 0;
            vector_output_0 = 0;
            vector_output_0[0] = out.s.y;
            vector_output_0[1] = out.s.x;
            vector_output_0[2] = in.s.x;
        }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

