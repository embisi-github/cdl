/*a Copyright
  
  This file 'vector_add.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/
constant integer width=16;

module vector_add( clock io_clock,
                     input bit io_reset,
                     input bit[width] vector_input_0,
                     input bit[width] vector_input_1,
                     output bit[width] vector_output_0,
                     output bit[width] vector_output_1 )
    "This module adds 1 to its vector output on every clock"
{
    default clock io_clock;
    default reset io_reset;

    clocked bit[width] vector_output_0 = 0;
    clocked bit[width] vector_output_1 = 0;

add_code:
    {
    vector_output_0 <= vector_output_0 + 1;
    }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

