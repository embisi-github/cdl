module reg( clock int_clock, input bit int_reset, input bit D, output bit Q )
{
    clocked clock rising int_clock reset active_high int_reset bit Q = 0;
    main_code "Main code":
        {
            Q <= D;
        }
}
