constant integer width=16;
typedef bit[width] value;
extern module adder( input value A, input value B, output value Z )
{
    timing comb input A, B;
    timing comb output Z;
}
module clocked_adder( clock int_clock,
                      input bit int_reset,
                      input value A,
                      input value B,
                      output value clocked_result
                     )
{
    net value result;
    clocked clock rising int_clock reset active_high int_reset value clocked_result = 0;

    instances "Adder instance":
        {
            adder add1( A<=A, B<=B, Z=>result );
        }
    registers "Register the result from the adder instance":
        {
            clocked_result <= result;
        }
}

