/*a Copyright
  
  This file 'vector_op_1.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/
constant integer width=16;
typedef bit[width] value;

module vector_op_1( clock io_clock,
                     input bit io_reset,
                     input value vector_input_0,
                     input value vector_input_1,
                     output value vector_output_0,
                     output value vector_output_1 )
    "This module sums uses bits of vector input 1 to decide whether to clear, add or subtract input 0 from output 0"
{
    default clock io_clock;
    default reset io_reset;

    clocked value vector_output_0 = 0;
    clocked value vector_output_1 = 0;
    comb value result;

generate_result:
    {
        result = vector_output_0;
        if (vector_input_1[0])
        {
            print("Clear result");
            result = 0;
        }
        if (vector_input_1[1])
        {
            print("Set result");
            result = vector_input_0;
        }
        if (vector_input_1[2])
        {
            print("Sum result and input");
            result = result + vector_input_0;
        }
        if (vector_input_1[3])
        {
            print("Subtract result and input");
            result = result - vector_input_0;
        }
    }
record_result:
    {
        vector_output_0 <= result;
    }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

