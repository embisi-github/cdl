/*a Copyright
  
  This file 'invert_chain.cdl' copyright Gavin J Stark 2003, 2004
  
  This program is free software; you can redistribute it and/or modify it under
  the terms of the GNU General Public License as published by the Free Software
  Foundation, version 2.0.
  
  This program is distributed in the hope that it will be useful,
  but WITHOUT ANY WARRANTY; without even implied warranty of MERCHANTABILITY
  or FITNESS FOR A PARTICULAR PURPOSE. See the GNU General Public License
  for more details.
*/
module invert_chain( input bit in_value,
                 output bit out_value_0,
                 output bit out_value_1,
                 output bit out_value_2,
                 output bit out_value_3,
                 output bit out_value_4,
                 output bit out_value_5,
                 output bit out_value_6,
                 output bit out_value_7
     )
    "This module implements a chain of inverters and outputs the results combinatorially"
{

invert_code:
    {
    out_value_4 = ~out_value_3;
    out_value_5 = ~out_value_4;

    out_value_7 = ~out_value_6;
    out_value_6 = ~out_value_5;

    out_value_0 = ~in_value;
    out_value_1 = ~out_value_0;
    out_value_2 = ~out_value_1;
    out_value_3 = ~out_value_2;
    }
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/

