constant integer fred=0;

constant bit bit=2;

constant a,b;

constant bit fjg=0

